`timescale 1ns / 1ps
module mips(clk, reset);
input clk;
input reset;

endmodule
